`ifndef CPU_DEFS_VH
`define CPU_DEFS_VH

`define ALU_CTRL_ADD  4'b0000
`define ALU_CTRL_SUB  4'b0001
`define ALU_CTRL_OR   4'b0010
`define ALU_CTRL_AND  4'b0011
`define ALU_CTRL_PASS 4'b0100

`define REG_RA        5'd31

`endif
